library ieee;
use ieee.std_logic_1164.all;

entity key_vector is
    port (
	index:		in     integer range 1 to 291;
	output:		out    std_logic_vector (1 to 64)
    );
end ;

architecture behave of key_vector is

    type vec_array is array (1 to 291) of std_logic_vector (1 to 64);

    constant vectors:	vec_array := (
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"0101010101010101",
	    x"8001010101010101",
	    x"4001010101010101",
	    x"2001010101010101",
	    x"1001010101010101",
	    x"0801010101010101",
	    x"0401010101010101",
	    x"0201010101010101",
	    x"0180010101010101",
	    x"0140010101010101",
	    x"0120010101010101",
	    x"0110010101010101",
	    x"0108010101010101",
	    x"0104010101010101",
	    x"0102010101010101",
	    x"0101800101010101",
	    x"0101400101010101",
	    x"0101200101010101",
	    x"0101100101010101",
	    x"0101080101010101",
	    x"0101040101010101",
	    x"0101020101010101",
	    x"0101018001010101",
	    x"0101014001010101",
	    x"0101012001010101",
	    x"0101011001010101",
	    x"0101010801010101",
	    x"0101010401010101",
	    x"0101010201010101",
	    x"0101010180010101",
	    x"0101010140010101",
	    x"0101010120010101",
	    x"0101010110010101",
	    x"0101010108010101",
	    x"0101010104010101",
	    x"0101010102010101",
	    x"0101010101800101",
	    x"0101010101400101",
	    x"0101010101200101",
	    x"0101010101100101",
	    x"0101010101080101",
	    x"0101010101040101",
	    x"0101010101020101",
	    x"0101010101018001",
	    x"0101010101014001",
	    x"0101010101012001",
	    x"0101010101011001",
	    x"0101010101010801",
	    x"0101010101010401",
	    x"0101010101010201",
	    x"0101010101010180",
	    x"0101010101010140",
	    x"0101010101010120",
	    x"0101010101010110",
	    x"0101010101010108",
	    x"0101010101010104",
	    x"0101010101010102",
	    x"8001010101010101",
	    x"4001010101010101",
	    x"2001010101010101",
	    x"1001010101010101",
	    x"0801010101010101",
	    x"0401010101010101",
	    x"0201010101010101",
	    x"0180010101010101",
	    x"0140010101010101",
	    x"0120010101010101",
	    x"0110010101010101",
	    x"0108010101010101",
	    x"0104010101010101",
	    x"0102010101010101",
	    x"0101800101010101",
	    x"0101400101010101",
	    x"0101200101010101",
	    x"0101100101010101",
	    x"0101080101010101",
	    x"0101040101010101",
	    x"0101020101010101",
	    x"0101018001010101",
	    x"0101014001010101",
	    x"0101012001010101",
	    x"0101011001010101",
	    x"0101010801010101",
	    x"0101010401010101",
	    x"0101010201010101",
	    x"0101010180010101",
	    x"0101010140010101",
	    x"0101010120010101",
	    x"0101010110010101",
	    x"0101010108010101",
	    x"0101010104010101",
	    x"0101010102010101",
	    x"0101010101800101",
	    x"0101010101400101",
	    x"0101010101200101",
	    x"0101010101100101",
	    x"0101010101080101",
	    x"0101010101040101",
	    x"0101010101020101",
	    x"0101010101018001",
	    x"0101010101014001",
	    x"0101010101012001",
	    x"0101010101011001",
	    x"0101010101010801",
	    x"0101010101010401",
	    x"0101010101010201",
	    x"0101010101010180",
	    x"0101010101010140",
	    x"0101010101010120",
	    x"0101010101010110",
	    x"0101010101010108",
	    x"0101010101010104",
	    x"0101010101010102",
	    x"1046913489980131",
	    x"1007103489988020",
	    x"10071034C8980120",
	    x"1046103489988020",
	    x"1086911519190101",
	    x"1086911519580101",
	    x"5107B01519580101",
	    x"1007B01519190101",
	    x"3107915498080101",
	    x"3107919498080101",
	    x"10079115B9080140",
	    x"3107911598080140",
	    x"1007D01589980101",
	    x"9107911589980101",
	    x"9107D01589190101",
	    x"1007D01598980120",
	    x"1007940498190101",
	    x"0107910491190401",
	    x"0107910491190101",
	    x"0107940491190401",
	    x"19079210981A0101",
	    x"1007911998190801",
	    x"10079119981A0801",
	    x"1007921098190101",
	    x"100791159819010B",
	    x"1004801598190101",
	    x"1004801598190102",
	    x"1004801598190108",
	    x"1002911498100104",
	    x"1002911598190104",
	    x"1002911598100201",
	    x"1002911698100101",
	    x"7CA110454A1A6E57",
	    x"0131D9619DC1376E",
	    x"07A1133E4A0B2686",
	    x"3849674C2602319E",
	    x"04B915BA43FEB5B6",
	    x"0113B970FD34F2CE",
	    x"0170F175468FB5E6",
	    x"43297FAD38E373FE",
	    x"07A7137045DA2A16",
	    x"04689104C2FD3B2F",
	    x"37D06BB516CB7546",
	    x"1F08260D1AC2465E",
	    x"584023641ABA6176",
	    x"025816164629B007",
	    x"49793EBC79B3258F",
	    x"4FB05E1515AB73A7",
	    x"49E95D6D4CA229BF",
	    x"018310DC409B26D6",
	    x"1C587F1C13924FEF"
	);
begin

    output <= vectors(index);

end behave;

