library ieee;
use ieee.std_logic_1164.all;

entity output_vector is
    port (
	index:		in     integer range 1 to 291;
	output:		out    std_logic_vector (1 to 64)
    );
end ;

architecture behave of output_vector is

    type vec_array is array (1 to 291) of std_logic_vector (1 to 64);

    constant vectors:	vec_array := (
	    x"8000000000000000",
	    x"4000000000000000",
	    x"2000000000000000",
	    x"1000000000000000",
	    x"0800000000000000",
	    x"0400000000000000",
	    x"0200000000000000",
	    x"0100000000000000",
	    x"0080000000000000",
	    x"0040000000000000",
	    x"0020000000000000",
	    x"0010000000000000",
	    x"0008000000000000",
	    x"0004000000000000",
	    x"0002000000000000",
	    x"0001000000000000",
	    x"0000800000000000",
	    x"0000400000000000",
	    x"0000200000000000",
	    x"0000100000000000",
	    x"0000080000000000",
	    x"0000040000000000",
	    x"0000020000000000",
	    x"0000010000000000",
	    x"0000008000000000",
	    x"0000004000000000",
	    x"0000002000000000",
	    x"0000001000000000",
	    x"0000000800000000",
	    x"0000000400000000",
	    x"0000000200000000",
	    x"0000000100000000",
	    x"0000000080000000",
	    x"0000000040000000",
	    x"0000000020000000",
	    x"0000000010000000",
	    x"0000000008000000",
	    x"0000000004000000",
	    x"0000000002000000",
	    x"0000000001000000",
	    x"0000000000800000",
	    x"0000000000400000",
	    x"0000000000200000",
	    x"0000000000100000",
	    x"0000000000080000",
	    x"0000000000040000",
	    x"0000000000020000",
	    x"0000000000010000",
	    x"0000000000008000",
	    x"0000000000004000",
	    x"0000000000002000",
	    x"0000000000001000",
	    x"0000000000000800",
	    x"0000000000000400",
	    x"0000000000000200",
	    x"0000000000000100",
	    x"0000000000000080",
	    x"0000000000000040",
	    x"0000000000000020",
	    x"0000000000000010",
	    x"0000000000000008",
	    x"0000000000000004",
	    x"0000000000000002",
	    x"0000000000000001",
	    x"95F8A5E5DD31D900",
	    x"DD7F121CA5015619",
	    x"2E8653104F3834EA",
	    x"4BD388FF6CD81D4F",
	    x"20B9E767B2FB1456",
	    x"55579380D77138EF",
	    x"6CC5DEFAAF04512F",
	    x"0D9F279BA5D87260",
	    x"D9031B0271BD5A0A",
	    x"424250B37C3DD951",
	    x"B8061B7ECD9A21E5",
	    x"F15D0F286B65BD28",
	    x"ADD0CC8D6E5DEBA1",
	    x"E6D5F82752AD63D1",
	    x"ECBFE3BD3F591A5E",
	    x"F356834379D165CD",
	    x"2B9F982F20037FA9",
	    x"889DE068A16F0BE6",
	    x"E19E275D846A1298",
	    x"329A8ED523D71AEC",
	    x"E7FCE22557D23C97",
	    x"12A9F5817FF2D65D",
	    x"A484C3AD38DC9C19",
	    x"FBE00A8A1EF8AD72",
	    x"750D079407521363",
	    x"64FEED9C724C2FAF",
	    x"F02B263B328E2B60",
	    x"9D64555A9A10B852",
	    x"D106FF0BED5255D7",
	    x"E1652C6B138C64A5",
	    x"E428581186EC8F46",
	    x"AEB5F5EDE22D1A36",
	    x"E943D7568AEC0C5C",
	    x"DF98C8276F54B04B",
	    x"B160E4680F6C696F",
	    x"FA0752B07D9C4AB8",
	    x"CA3A2B036DBC8502",
	    x"5E0905517BB59BCF",
	    x"814EEB3B91D90726",
	    x"4D49DB1532919C9F",
	    x"25EB5FC3F8CF0621",
	    x"AB6A20C0620D1C6F",
	    x"79E90DBC98F92CCA",
	    x"866ECEDD8072BB0E",
	    x"8B54536F2F3E64A8",
	    x"EA51D3975595B86B",
	    x"CAFFC6AC4542DE31",
	    x"8DD45A2DDF90796C",
	    x"1029D55E880EC2D0",
	    x"5D86CB23639DBEA9",
	    x"1D1CA853AE7C0C5F",
	    x"CE332329248F3228",
	    x"8405D1ABE24FB942",
	    x"E643D78090CA4207",
	    x"48221B9937748A23",
	    x"DD7C0BBD61FAFD54",
	    x"2FBC291A570DB5C4",
	    x"E07C30D7E4E26E12",
	    x"0953E2258E8E90A1",
	    x"5B711BC4CEEBF2EE",
	    x"CC083F1E6D9E85F6",
	    x"D2FD8867D50D2DFE",
	    x"06E7EA22CE92708F",
	    x"166B40B44ABA4BD6",
	    x"95A8D72813DAA94D",
	    x"0EEC1487DD8C26D5",
	    x"7AD16FFB79C45926",
	    x"D3746294CA6A6CF3",
	    x"809F5F873C1FD761",
	    x"C02FAFFEC989D1FC",
	    x"4615AA1D33E72F10",
	    x"2055123350C00858",
	    x"DF3B99D6577397C8",
	    x"31FE17369B5288C9",
	    x"DFDD3CC64DAE1642",
	    x"178C83CE2B399D94",
	    x"50F636324A9B7F80",
	    x"A8468EE3BC18F06D",
	    x"A2DC9E92FD3CDE92",
	    x"CAC09F797D031287",
	    x"90BA680B22AEB525",
	    x"CE7A24F350E280B6",
	    x"882BFF0AA01A0B87",
	    x"25610288924511C2",
	    x"C71516C29C75D170",
	    x"5199C29A52C9F059",
	    x"C22F0A294A71F29F",
	    x"EE371483714C02EA",
	    x"A81FBD448F9E522F",
	    x"4F644C92E192DFED",
	    x"1AFA9A66A6DF92AE",
	    x"B3C1CC715CB879D8",
	    x"19D032E64AB0BD8B",
	    x"3CFAA7A7DC8720DC",
	    x"B7265F7F447AC6F3",
	    x"9DB73B3C0D163F54",
	    x"8181B65BABF4A975",
	    x"93C9B64042EAA240",
	    x"5570530829705592",
	    x"8638809E878787A0",
	    x"41B9A79AF79AC208",
	    x"7A9BE42F2009A892",
	    x"29038D56BA6D2745",
	    x"5495C6ABF1E5DF51",
	    x"AE13DBD561488933",
	    x"024D1FFA8904E389",
	    x"D1399712F99BF02E",
	    x"14C1D7C1CFFEC79E",
	    x"1DE5279DAE3BED6F",
	    x"E941A33F85501303",
	    x"DA99DBBC9A03F379",
	    x"B7FC92F91D8E92E9",
	    x"AE8E5CAA3CA04E85",
	    x"9CC62DF43B6EED74",
	    x"D863DBB5C59A91A0",
	    x"A1AB2190545B91D7",
	    x"0875041E64C570F7",
	    x"5A594528BEBEF1CC",
	    x"FCDB3291DE21F0C0",
	    x"869EFD7F9F265A09",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"0000000000000000",
	    x"88D55E54F54C97B4",
	    x"0C0CC00C83EA48FD",
	    x"83BC8EF3A6570183",
	    x"DF725DCAD94EA2E9",
	    x"E652B53B550BE8B0",
	    x"AF527120C485CBB0",
	    x"0F04CE393DB926D5",
	    x"C9F00FFC74079067",
	    x"7CFD82A593252B4E",
	    x"CB49A2F9E91363E3",
	    x"00B588BE70D23F56",
	    x"406A9A6AB43399AE",
	    x"6CB773611DCA9ADA",
	    x"67FD21C17DBB5D70",
	    x"9592CB4110430787",
	    x"A6B7FF68A318DDD3",
	    x"4D102196C914CA16",
	    x"2DFA9F4573594965",
	    x"B46604816C0E0774",
	    x"6E7E6221A4F34E87",
	    x"AA85E74643233199",
	    x"2E5A19DB4D1962D6",
	    x"23A866A809D30894",
	    x"D812D961F017D320",
	    x"055605816E58608F",
	    x"ABD88E8B1B7716F1",
	    x"537AC95BE69DA1E1",
	    x"AED0F6AE3C25CDD8",
	    x"B3E35A5EE53E7B8D",
	    x"61C79C71921A2EF8",
	    x"E2F5728F0995013C",
	    x"1AEAC39A61F0A464",
	    x"690F5B0D9A26939B",
	    x"7A389D10354BD271",
	    x"868EBB51CAB4599A",
	    x"7178876E01F19B2A",
	    x"AF37FB421F8C4095",
	    x"86A560F10EC6D85B",
	    x"0CD3DA020021DC09",
	    x"EA676B2CB7DB2B7A",
	    x"DFD64A815CAF1A0F",
	    x"5C513C9C4886C088",
	    x"0A2AEEAE3FF4AB77",
	    x"EF1BF03E5DFA575A",
	    x"88BF0DB6D70DEE56",
	    x"A1F9915541020B56",
	    x"6FBF1CAFCFFD0556",
	    x"2F22E49BAB7CA1AC",
	    x"5A6B612CC26CCE4A",
	    x"5F4C038ED12B2E41",
	    x"63FAC0D034D9F793"
	);
begin

    output <= vectors(index);

end behave;

