library ieee;
use ieee.std_logic_1164.all;

entity encrypt_vector is
    port (
	index:		in     integer range 1 to 291;
	output:		out    std_logic
    );
end ;

architecture behave of encrypt_vector is

    constant bit_array:	std_logic_vector(1 to 291) := (
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0',
	    '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
	    '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
	    '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1',
	    '1','1','1'
	);
    begin

    output <= bit_array(index);

end behave;

